`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/01/2025 05:13:43 PM
// Design Name: 
// Module Name: imgen
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
//==============================================================
// Immediate Generator for RISC-V Processor
//==============================================================
module imgen (
    input  [31:0] instr,      // 32-bit instruction
    output reg [31:0] imm_out // 32-bit immediate output
);

    wire [6:0] opcode = instr[6:0];

    always @(*) begin
        case (opcode)
            7'b0000011, // I-type (LW)
            7'b0010011, // I-type (ADDI)
            7'b1100111: // I-type (JALR)
                imm_out = {{20{instr[31]}}, instr[31:20]};

            7'b0100011: // S-type (SW)
                imm_out = {{20{instr[31]}}, instr[31:25], instr[11:7]};

            7'b1100011: // B-type (BEQ)
                imm_out = {{19{instr[31]}}, instr[31], instr[7],
                           instr[30:25], instr[11:8], 1'b0};

            7'b0110111, // U-type (LUI)
            7'b0010111: // U-type (AUIPC)
                imm_out = {instr[31:12], 12'b0};

            7'b1101111: // J-type (JAL)
                imm_out = {{11{instr[31]}}, instr[31],
                           instr[19:12], instr[20], instr[30:21], 1'b0};

            default:
                imm_out = 32'b0;
        endcase
    end
endmodule

